
module SignedMultiplier_ShiftAdd_AxB(
	);
	
	
endmodule