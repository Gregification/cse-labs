/**
	cse3341, digital logic 2, lab 5
	George Boone
	1002055713

	modular exponent subtractor
	this module is not part of the logic, it only serves to demo it
*/

module lab5(
		// standard in. i got tired of the assignment editor, see immideatly after wire decelerations for assignments
		input [9:0] DEVBOARD_SWS,
		input [1:0] DEVBOARD_BTN,
		output[9:0] DEVBOARD_RLEDS,	
		output[47:0]DEBBOARD_SEGS,
		input [3:0] HEXBOARD_BTN,	
		output[3:0] HEXBOARD_CAT,
		output[6:0] HEXBOARD_SEGS
	);
	
	
//------------------------------------------------------------------------------
// 	INPUT ASSIGMENTS  \ EXTERNAL WIRING
//------------------------------------------------------------------------------

	wire [7:0] _input_value;
	
//------------------------------------------------------------------------------
// 	INTERNAL WIRING
//------------------------------------------------------------------------------	


//------------------------------------------------------------------------------
// 	MODULES
//------------------------------------------------------------------------------	
	
endmodule
