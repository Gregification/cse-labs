/**
cse3341, digital logic 2, lab 4
George Boone
1002055713
*/

module lab4(
	);
	
endmodule
