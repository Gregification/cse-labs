
module lab4(
	);
	
endmodule;
